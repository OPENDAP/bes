netcdf fnoc_hacked {
dimensions:
	lat = 17 ;
	lon = 21 ;
variables:
	short u(lat, lon) ;
		u:units = "meter per second" ;
		u:long_name = "Vector wind eastward component" ;
		u:missing_value = "-32767" ;
		u:scale_factor = "0.005" ;
	short v(lat, lon) ;
		v:units = "meter per second" ;
		v:long_name = "Vector wind northward component" ;
		v:missing_value = "-32767" ;
		v:scale_factor = "0.005" ;
	float lat(lat) ;
		lat:units = "degree North" ;
	float lon(lon) ;
		lon:units = "degree East" ;

// global attributes:
		:base_time = "88- 10-00:00:00" ;
		:title = " FNOC UV wind components from 1988- 10 to 1988- 13." ;
data:

 u =
  -1728, -2449, -3099, -3585, -3254, -2406, -1252, 662, 2483, 2910, 2819, 
    2946, 2745, 2734, 2931, 2601, 2139, 1845, 1754, 1897, 1854,
  -1686, -1985, -2508, -3397, -3501, -3268, -2700, -705, 1834, 2728, 2484, 
    2465, 2531, 2591, 2514, 2200, 1934, 1677, 1401, 1202, 1084,
  -223, -864, -864, -1152, -1427, -1717, -1992, -1211, 791, 2235, 2558, 2770, 
    2961, 2663, 2131, 1959, 2035, 2053, 1732, 926, 581,
  1924, 1664, 1555, 1551, 1190, 430, -459, -453, 914, 2055, 2526, 2916, 2761, 
    1955, 1418, 1509, 1645, 1720, 1510, 739, 318,
  2869, 3660, 3561, 3069, 2378, 1453, 601, 479, 953, 1237, 1494, 1700, 1436, 
    751, 358, 732, 1067, 922, 701, 484, 166,
  2012, 2885, 3172, 2734, 2141, 1453, 795, 420, -98, -415, -37, 108, -104, 
    -313, -609, -225, 559, 508, 144, 128, -57,
  685, 1311, 1566, 1458, 1174, 762, 327, -113, -779, -1281, -1168, -968, 
    -932, -1048, -1344, -1051, -235, 72, -14, -6, -83,
  -135, 336, 408, 261, -1, -305, -509, -664, -932, -1326, -1734, -1680, 
    -1197, -1260, -1784, -1724, -1132, -545, -169, -26, 92,
  -628, -593, -482, -575, -792, -1064, -1290, -1280, -1125, -1202, -1598, 
    -1676, -1340, -1307, -1652, -1748, -1393, -896, -534, -363, -175,
  -903, -1244, -1158, -1036, -1219, -1432, -1556, -1551, -1223, -1041, -1074, 
    -1040, -1194, -1380, -1351, -1211, -916, -749, -956, -1132, -1125,
  -1247, -1435, -1261, -1147, -1445, -1657, -1641, -1599, -1298, -1042, -946, 
    -630, -512, -1018, -1489, -1185, -483, -401, -1168, -1888, -2185,
  -1873, -1883, -1557, -1411, -1469, -1584, -1648, -1599, -1362, -1119, 
    -1068, -760, -282, -690, -1633, -1489, -569, -324, -906, -1711, -2371,
  -2116, -2318, -2171, -1834, -1610, -1576, -1672, -1547, -1307, -1238, 
    -1113, -936, -745, -782, -1320, -1385, -635, -48, -131, -907, -1877,
  -2055, -2123, -2049, -1781, -1842, -2019, -2132, -1775, -1288, -1227, 
    -1023, -787, -848, -845, -1010, -1162, -522, 403, 488, -509, -1602,
  -2087, -1807, -1623, -1734, -1891, -2086, -2257, -1897, -1349, -1079, -811, 
    -698, -1040, -1163, -933, -944, -617, 193, 388, -413, -1269,
  -1942, -1670, -1472, -1896, -1915, -1669, -1709, -1607, -1319, -1140, -959, 
    -911, -1290, -1252, -467, -281, -597, -429, -251, -484, -749,
  -1661, -1294, -934, -1328, -1643, -1426, -1321, -1400, -1250, -1130, -1209, 
    -1096, -929, -669, 42, 212, -485, -892, -865, -605, -303;

 v =
  -2067, -2025, -668, 603, 1419, 2261, 2410, 1566, 429, -286, -475, -838, 
    -1354, -1373, -969, -524, -28, 452, 640, 618, 595,
  -3100, -3037, -999, 1124, 2528, 3511, 3779, 2626, 695, -340, -579, -780, 
    -833, -915, -1144, -982, -279, 344, 510, 291, -2,
  -3139, -3255, -750, 1608, 2788, 3856, 4321, 3137, 1477, 692, 200, -123, 
    -252, -919, -1623, -1334, -385, 432, 708, 201, -328,
  -2858, -2657, -155, 2000, 3020, 4009, 4239, 3193, 1562, 483, 265, 105, 
    -456, -1483, -2014, -1368, -373, 471, 740, 224, -139,
  -1812, -1465, 362, 2554, 3907, 4324, 4030, 3236, 1379, -376, -547, -564, 
    -1144, -1751, -1939, -1405, -651, 2, 266, 141, 63,
  -511, -288, 1165, 3002, 3738, 3543, 3070, 2283, 1194, 17, -798, -1211, 
    -1345, -1348, -1471, -1617, -1497, -747, 12, 114, -40,
  335, 570, 1698, 2684, 2511, 1891, 1384, 698, 337, 130, -635, -1090, -855, 
    -953, -1401, -1825, -1995, -1011, 201, 235, -16,
  776, 901, 1179, 1530, 1528, 981, 331, -209, -640, -706, -731, -764, -539, 
    -721, -1419, -1868, -1785, -991, 46, 353, 231,
  891, 570, 231, 619, 1169, 874, 189, -370, -982, -1198, -792, -517, -463, 
    -403, -898, -1505, -1338, -781, -175, 256, 299,
  614, 44, -232, 314, 816, 410, -83, -356, -857, -1158, -747, -256, -245, 
    -457, -875, -1137, -734, -198, -35, 9, 108,
  97, -206, -208, -51, -32, -459, -687, -531, -649, -982, -833, -270, -257, 
    -1092, -1680, -1157, -259, 110, 135, 110, -69,
  -304, -342, -292, -421, -627, -802, -856, -747, -740, -895, -864, -562, 
    -560, -1393, -2086, -1354, -320, -125, 115, 348, -153,
  -425, -325, -399, -606, -713, -679, -730, -892, -989, -915, -738, -763, 
    -865, -1108, -1557, -1276, -544, -306, -102, 27, -407,
  -123, -68, -262, -579, -651, -751, -830, -922, -1085, -1004, -710, -734, 
    -994, -997, -821, -604, -317, -178, -273, -500, -811,
  145, -90, -282, -449, -555, -653, -687, -823, -1017, -963, -775, -702, 
    -855, -934, -623, -338, -240, -204, -356, -635, -917,
  110, -224, -374, -422, -517, -309, -347, -640, -640, -711, -782, -620, 
    -663, -792, -756, -729, -635, -524, -477, -414, -527,
  345, 96, -107, -149, -220, -333, -437, -346, -397, -768, -584, -185, -629, 
    -1203, -1068, -628, -493, -719, -646, 19, 356;

 lat = 50, 47.5, 45, 42.5, 40, 37.5, 35, 32.5, 30, 27.5, 25, 22.5, 20, 17.5, 
    15, 12.5, 10 ;

 lon = -60, -57.5, -55, -52.5, -50, -47.5, -45, -42.5, -40, -37.5, -35, 
    -32.5, -30, -27.5, -25, -22.5, -20, -17.5, -15, -12.5, -10 ;
}

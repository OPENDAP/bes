netcdf ref_tst_compounds3 {
types:
  compound cmp1 {
    short i ;
    int j ;
  }; // cmp1
  compound cmp2 {
    float x ;
    double y ;
  }; // cmp2
  compound cmp3 {
    cmp1 xx ;
    cmp2 yy ;
  }; // cmp3

variables:
	cmp3 phony_compound_var ;
        phony_compound_var:desc="A scalar nested compound dataset";
data:

 phony_compound_var = 
    {{20000, 300000}, {100000, -100000.028899567}};
}

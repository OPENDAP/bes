netcdf ref_tst_compounds5 {
types:
  compound cmp1 {
    short i ;
    int j ;
  }; // cmp1
  compound cmp2 {
    float x ;
    double y(3, 2) ;
  }; // cmp2
  compound cmp3 {
    cmp1 xx ;
    cmp2 yy ;
  }; // cmp3
dimensions:
	phony_dim = 2 ;
variables:
	cmp3 phony_compound_var(phony_dim) ;
data:

 phony_compound_var =
     {{20000, 300000}, {100000, {-100000.028899567, -200000, -300000, -400000, -500000, 3.1415926}}},
     {{20000, 300000}, {100000, {-100000.028899567, -100000, -100000, -100000, -100000, -100000}}};
}

netcdf group_mlls{
dimensions:
        lat = 2 ;
        lon = 3 ;
variables:
        float lat(lat);
              lat:units = "degrees_north";
        float lon(lon);
              lon:units = "degrees_east";
        float pres1(lat,lon);
              pres1:units = "hPa";
data:
        lat = 2,4;
        lon = -10,-5,0;
        pres1 =
          900,902,904,
          901,903,905;
group: g1 {
 dimensions:
       dim1 = 4;
       dim2 = 6;
 variables:
   int dim1(dim1);
   int dim2(dim2);
   float lat1(dim1,dim2);
         lat1:units = "degrees_north";
   float lon1(dim1,dim2);
         lon1:units = "degrees_east";
   float pres2(dim1,dim2);
         pres2:units = "hPa";
 data:
       dim1 = 1,2,3,4;
       dim2 = 1,2,3,4,5,6;
       lat1 = 2,2.5,3,3.5,5,6,
              2.1,2.6,3.1,3.6,5.1,6.1,
              2.4,2.9,3.4,3.9,5.4,6.4,
              2.8,3.3,3.8,4.3,5.8,6.8;
       lon1 = -10,-8,-6,-4,3,4,
              -9,-7,-5,-3,4,5,
              -6,-4,-1,0,7,8,
              -4,-2,1,2,9,10;
       pres2 = 800,810,820,830,840,850,
               801,811,821,831,841,851,
               802,812,822,832,842,852,
               803,813,823,833,843,853;
 }
group: g2 {
 dimensions:
       dim1 = 2;
       dim2 = 3;
 variables:
   float lat1(dim1,dim2);
         lat1:units = "degrees_north";
   float lon1(dim1,dim2);
         lon1:units = "degrees_east";
   float temp1(dim1,dim2);
         temp1:units = "K";
 data:
       lat1 = 2,3,5,
              2.8,3.8,5.8;
       lon1 = -10,-6,3,
              -6,-1,7;
       temp1 = 271,272,273,
               270,271,272;
}
group: g3 {
 dimensions:
       dim1 = 2;
       dim2 = 3;
 variables:
   float latitude(dim1,dim2);
   float longitude(dim1,dim2);
   float temp2(dim1,dim2);
         temp2:units = "K";
 data:
       latitude = -2,-3,-5,
              -2.1,-3.1,-5.1;
       longitude = 10,6,3,
              16,20,27;
       temp2 = 261,262,263,
               260,261,262;
}
}

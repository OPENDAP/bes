netcdf comp_complex_scalar {
types:
  compound cmp1 {
    short i ;
    int j ;
  }; // cmp1
  compound cmp2 {
    float f;
    cmp1 x ;
    double y(2) ;
  }; // cmp2
  compound cmp3 {
    cmp2 yy(5) ;
  }; // cmp3

variables:
	cmp3 phony_compound_var;
data:
 phony_compound_var = 
    {{{1.1, {1, 20000}, {-100000.285657, 3.1415926}},
      {2.2, {2, 40000}, {-200000.285657, 4.1415926}},
      {3.3, {3, 60000}, {-300000.285657, 5.1415926}},
      {5.5, {4, 80000}, {-400000.285657, 6.1415926}},
      {6.6, {5, 100000},{-500000.285657, 7.1415926}}}}; 
}


netcdf test {

dimensions:
	nodes = 9 ;

variables:
	float X(nodes) ;

data:
 
 X = -1.0, 0.0, 1.0, 1.5,  1.0,  0.0, -1.0, -1.5, 0.0 ;

}

netcdf compound_array_complex_more {
types:
  compound cmp1 {
    short i ;
    int j ;
  }; // cmp1
  compound cmp2 {
    cmp1 x ;
    double y(3) ;
  }; // cmp2
  compound cmp3 {
    cmp2 yy(3) ;
  }; // cmp3
dimensions:
   n=4;

variables:
	cmp3 phony_compound_var(n);
data:

 phony_compound_var = 
    
    {{{{1, 100000}, {100000.285657, 100.1, 1.1415926}},
      {{2,200000},  {200000.151617,200.2,273.15}},
      {{-1, -100000}, {-100000.285657, -100.1,-1.1415926}}}}, 
    {{{{3, 300000}, {300000.285657, 300.3, 3.1415926}},
      {{4,400000},  {400000.151617,400.4,473.15}},
      {{-2, -200000}, {-200000.285657, -200.2,-2.1415926}}}}, 
    {{{{5, 500000}, {500000.285657, 500.5, 5.1415926}},
      {{6,600000},  {600000.151617,600.6,673.15}},
      {{-3, -300000}, {-300000.285657, -300.3,-3.1415926}}}}, 
    {{{{7, 700000}, {700000.275657, 700.7, 7.1415926}},
      {{8,800000},  {800000.151617,800.8,873.15}},
      {{-4, -400000}, {-400000.285657, -400.4,-4.1415926}}}}; 
}

netcdf t_group {
dimensions:
        dim1 = 2 ;
        dim2 = 3 ;
 group: g1 {
  variables:
   float d1(dim1,dim2);
   d1:coordinates = "/g2/c1 /g2/c2";
   float d2(dim1,dim2);
   d2:coordinates = "g2/c3 g2/c4";
  data:
       d1 = 0.5,1.5,2.5,3.5,4.5,5.5;
       d2 = 6.5,7.5,8.5,9.5,10.5,11.5;
 }
 group: g2 {
   variables:
    int c1(dim1,dim2);
    int c2(dim1,dim2);
    int c3(dim1,dim2);
    int c4(dim1,dim2);
   data:
       c1 = 1,2,3,4,5,6;
       c2 = 2,3,4,5,6,7;
       c3 = 3,4,5,6,7,8;
       c4 = 4,5,6,7,8,9;
 }
}

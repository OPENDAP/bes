netcdf group_mlls_nocvs{
dimensions:
        dimr0 = 2 ;
        dimr1 = 3 ;
variables:
        float lat1(dimr0,dimr1);
              lat1:units = "degrees_north";
        float lon1(dimr0,dimr1);
              lon1:units = "degrees_east";
        float lat2(dimr0,dimr1);
              lat2:units = "degrees_north";
        float lon2(dimr0,dimr1);
              lon2:units ="degrees_east";
        float pres1(dimr0,dimr1);
              pres1:units = "hPa";
              pres1:coordinates="/lat1 /lon1";
        float pres2(dimr0,dimr1);
              pres2:units = "hPa";

data:
        lat1 = 1,2,3,4,5,6;
        lon1 = 2,4,6,8,10,12;
        lat2 = -1,-2,-3,-4,-5,-6;
        lon2 = -2,-4,-6,-8,-10,-12;
        pres1 =
          900,902,904,
          901,903,905;
        pres2 =
          1000,1001,1002,
          1003,1004,1005;
group: g1 {
 dimensions:
       dim1 = 2;
       dim2 = 3;
 variables:
   int dim1(dim1);
   int dim2(dim2);
   float lat1(dim1,dim2);
         lat1:units = "degrees_north";
   float lat2(dim1,dim2);
         lat2:units = "degrees_north";
   float lon1(dim1,dim2);
         lon1:units = "degrees_east";
   float pres2(dim1,dim2);
         pres2:units = "hPa";
 data:
       dim1 = 1,2;
       dim2 = 1,2,3;
       lat1 = 2,2.5,3,3.5,5,6;
       lat2 = 4,4.5,6,6.5,7,8;
       lon1 = -10,-8,-6,-4,3,4;
       pres2 = 800,810,820,830,840,850;
 }
group: g2 {
 dimensions:
       dim1 = 2;
       dim2 = 3;
 variables:
   float lon1(dim1,dim2);
         lon1:units = "degrees_east";
   float temp1(dim1,dim2);
         temp1:units = "K";
 data:
       lon1 = -10,-6,3,
              -6,-1,7;
       temp1 = 271,272,273,
               270,271,272;
}
group: g3 {
 dimensions:
       dim1 = 2;
       dim2 = 3;
 variables:
   float lat1(dim1,dim2);
         lat1:units="degrees_east";
   float lon1(dim1,dim2);
         lon1:units="degrees_north";
   float lat2(dim1,dim2);
         lat2:units="degrees_east";
   float lon2(dim1,dim2);
         lon2:units="degrees_north";
  float temp1(dim1,dim2);
         temp1:units = "K";
         temp1:coordinates="/g3/lat1 /g3/lon1";
  float temp2(dim1,dim2);
         temp2:units = "K";
data:
       lat1 = -2,-3,-5,
              -2.1,-3.1,-5.1;
       lon1 = 10,6,3,
              16,20,27;
        lat2 = -2,-3,-5,
              -2.1,-3.1,-5.1;
       lon2 = 10,6,3,
              16,20,27;
      temp1 = 271,272,273,274,275,276;
      temp2 = 261,262,263,
               260,261,262;
}
}

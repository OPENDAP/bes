netcdf group_mlls_sdim{
dimensions:
        dim0 = 4 ;
        dim1 = 3;
variables:
        float latitude(dim0,dim1);
        float longitude(dim0,dim1);
data:
       latitude = 80,81,82,
                  81,82,83,
                  82,83,84,
                  83,84,85;
       longitude = 120,121,122,
                   121,122,123,
                   122,123,124,
                   123,124,125;
                  
group: g1 {
 dimensions:
       dim1 = 6;
 variables:
   int dim1(dim1);
   float lat1(dim0,dim1);
         lat1:units = "degrees_north";
   float lon1(dim0,dim1);
         lon1:units = "degrees_east";
   float pres2(dim0,dim1);
         pres2:units = "hPa";
 data:
       dim1 = 1,2,3,4,5,6;
       lat1 = 2,2.5,3,3.5,5,6,
              2.1,2.6,3.1,3.6,5.1,6.1,
              2.4,2.9,3.4,3.9,5.4,6.4,
              2.8,3.3,3.8,4.3,5.8,6.8;
       lon1 = -10,-8,-6,-4,3,4,
              -9,-7,-5,-3,4,5,
              -6,-4,-1,0,7,8,
              -4,-2,1,2,9,10;
       pres2 = 800,810,820,830,840,850,
               801,811,821,831,841,851,
               802,812,822,832,842,852,
               803,813,823,833,843,853;
 }
group: g2 {
 dimensions:
       dim1 = 2;
 variables:
   float lat1(dim1,dim0);
         lat1:units = "degrees_north";
   float lon1(dim1,dim0);
         lon1:units = "degrees_east";
   float temp1(dim1,dim0);
         temp1:units = "K";
 data:
       lat1 = 2,3,5,6,
              2.8,3.8,5.8,6.8;
       lon1 = -10,-6,3,3.1,
              -6,-1,7,8;
       temp1 = 271,272,273,274,
               270,271,272,273;
}
group: g3 {
 variables:
   float temp2(dim0,dim1);
         temp2:units = "K";
 data:
       temp2 = 280,281,282,
               281,282,283,
               282,283,284,
               283,284,285;
}
}
